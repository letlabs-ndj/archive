LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY bcd IS PORT (
	I: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	S: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	N: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	Segs: OUT std_logic_vector (1 TO 7));
END bcd;

ARCHITECTURE Behavioral OF bcd IS
BEGIN
	PROCESS(I,S,N)
	BEGIN
		CASE I IS
		WHEN "00000" => Segs <= "11110011001100000000";
		WHEN "00001" => Segs <= "10011111101100000000";
		WHEN "00010" => Segs <= "11001111000000000000";
		WHEN "00011" => Segs <= "10011111000000000000";
		WHEN "00100" => Segs <= "11001111001100000000";
		WHEN "00101" => Segs <= "11000011001100000000";
		WHEN "00110" => Segs <= "11011111000100000000";
		WHEN "00111" => Segs <= "00110011001100000000";
		WHEN "01000" => Segs <= "00000000110000000000";
		WHEN "01001" => Segs <= "00111110000000000000";
		WHEN "01010" => Segs <= "00000000110000000000";
		WHEN "01011" => Segs <= "00001111000000000000";
		WHEN "01100" => Segs <= "00110011000010100000";
		WHEN "01101" => Segs <= "00110011000011000000";
		WHEN "01110" => Segs <= "11111111000000000000";
		WHEN "01111" => Segs <= "11100011001100000000";
		WHEN "10000" => Segs <= "11111111000001000000";
		WHEN "10001" => Segs <= "11100011000010100000";
		WHEN "10010" => Segs <= "11011101001100000000";
		WHEN "10011" => Segs <= "11000000110000000000";
		WHEN "10100" => Segs <= "00111111000000000000";
		WHEN "10101" => Segs <= "00100001000000000000";
		WHEN "10110" => Segs <= "00110011000001010000";
		WHEN "10111" => Segs <= "00000000000011110000";
		WHEN "11000" => Segs <= "00000000010010100000";
		WHEN OTHERS => Segs <= "11001100000000110000";
		END CASE;
	END PROCESS;
END Behavioral;
